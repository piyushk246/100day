module johnson();

endmodule
